`ifndef REG_SEQUENCER_SVH
`define REG_SEQUENCER_SVH

//-----------------------------------------------------------------------------
// Class: reg_sequencer
// Description: UVM sequencer for register transactions
//-----------------------------------------------------------------------------

typedef uvm_sequencer #(reg_item) reg_sequencer;

`endif
